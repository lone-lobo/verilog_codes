module ();
input ;
output ;

parameters ;

case ()
  
  
  default:begin
  end
  

endmodule
